// file pipelineIF_ID_Register.v

module pipelineIF_ID_Register(
	input wire clock,
	input wire [31:0] instr);